module seven_segment_decoder (
    input logic [3:0] D,        // 4-bit binary input representing hexadecimal digit
    input logic RBI,            // Ripple Blanking Input
    output logic [6:0] seg,     // 7-segment outputs: seg[6] = a, ..., seg[0] = g (active low)
    output logic RBO            // Ripple Blanking Output
);
    logic zero; // flag for input D = 0

    always_comb begin
        // Default case: inactive segments (all off = all high, since active low)
        seg = 7'b1111111;
        zero = (D == 4'd0);

        case (D)
            4'h0: seg = 7'b1111110;
            4'h1: seg = 7'b0110000;
            4'h2: seg = 7'b1101101;
            4'h3: seg = 7'b1111001;
            4'h4: seg = 7'b0110011;
            4'h5: seg = 7'b1011011;
            4'h6: seg = 7'b1011111;
            4'h7: seg = 7'b1110000;
            4'h8: seg = 7'b1111111;
            4'h9: seg = 7'b1110011;
            4'hA: seg = 7'b1110111;
            4'hB: seg = 7'b0011111;
            4'hC: seg = 7'b1001110;
            4'hD: seg = 7'b0111101;
            4'hE: seg = 7'b1001111;
            4'hF: seg = 7'b1000111;
        endcase

        // Ripple blanking logic: suppress 0 if RBI = 0
        if (zero && !RBI)
            seg = 7'b1111111; // Blank the display

        // Set RBO: should propagate 0 suppression
        RBO = zero && !RBI;
    end
endmodule